//////////////////////////////////////////////////////////////
////////////////       Transaction Class       ///////////////
//////////////////////////////////////////////////////////////
class Transaction #(
    
                    parameter Data_Width = 32,
					parameter Addr_Width = 5 
                        
                    );

/*

    Description:    Defines the pin level activity generated by agent (to drive to DUT through the driver) or 
                    the activity has to be observed by agent 

*/

         
	rand  bit			     		 Wr_En    ;
	rand  bit			     		 Rd_En    ;
	rand  bit 	[Data_Width - 1 : 0] Data_in  ;
	randc bit 	[Addr_Width - 1 : 0] Address  ;
	      bit   [Data_Width - 1 : 0] Data_out ;
	      bit   		             Valid_out;
		  bit 						 cnt	  ;
		 
	constraint value_A {Address inside {['d0:'d31]};}
	constraint wr_rd_C { Wr_En != Rd_En; };
    
    function new ();
        
    endfunction

    function void print (string tag="");

        $display("T = %0t [%s] \t Address = %0d \t Wr_En = %d \t Data_in = %0h \t Rd_En = %0d \t Data_out = %0h \n", $time, tag, Address, Wr_En, Data_in, Rd_En, Data_out);
        $display(" --------------------------------------------------------- \n");

    endfunction  
  
endclass //Transaction
