////////////////////////////////////////////////////////////
// Author	: Mahmoud Magdi 
// Date  	: 11 - Nov. - 2023
// Version 	: Stable
////////////////////////////////////////////////////////////



`define DRIV_IF mem_vif.DRIVER.Driver_cb					// `DRIV_IF will point to mem_vif.DRIVER.Driver_cb which is in the virtual interface
`define MONT_IF mem_vif.MONITOR.Monitor_cb

//////////////////////////////////////////////////////////////
////////////////       Transaction Class       ///////////////
//////////////////////////////////////////////////////////////
class Transaction #(
    
                    parameter Data_Width = 32,
					parameter Addr_Width = 5 
                        
                    );

/*

    Description:    Defines the pin level activity generated by agent (to drive to DUT through the driver) or 
                    the activity has to be observed by agent 

*/

         
	rand  bit			     		 Wr_En    ;
	rand  bit			     		 Rd_En    ;
	rand  bit 	[Data_Width - 1 : 0] Data_in  ;
	randc bit 	[Addr_Width - 1 : 0] Address  ;
	      bit   [Data_Width - 1 : 0] Data_out ;
	      bit   		             Valid_out;
		  bit 						 cnt	  ;
		 
	constraint value_A {Address inside {['d0:'d31]};}
	constraint wr_rd_C { Wr_En != Rd_En; };
    
    function new ();
        
    endfunction

    function void print (string tag="");

        $display("T = %0t [%s] \t Address = %0d \t Wr_En = %d \t Data_in = %0h \t Rd_En = %0d \t Data_out = %0h \n", $time, tag, Address, Wr_En, Data_in, Rd_En, Data_out);
        $display(" --------------------------------------------------------- \n");

    endfunction  
  
endclass //Transaction






//////////////////////////////////////////////////////////////
////////////////        Sequencer Class        ///////////////
//////////////////////////////////////////////////////////////
class Sequencer;

	rand Transaction #(32,5)trn;
	
	
	// Creating a Mailbox is used to send the randomized transaction to Driver
	mailbox mbox;
    
	// Adding a variable to control the number of random packets to be created
	int repeat_count;
	
	
	//  Adding an event to indicate the completion of the generation process, 
	//  the event will be triggered on the completion of the Generation process.
	event completed;
	
	
	// Constructor
	function new(mailbox mbox, event completed);			
        
		// getting the mailbox handle from env
		this.mbox   = mbox;
		this.completed = completed;
		
    endfunction //new()

	

	// Main task that creates and randomize the stimulus and puts into the mailbox
    task stimulus ();
	
		repeat(repeat_count)
		begin
		
			trn = new();
			// trn.randomize();
			if (!trn.randomize ()) $fatal("Gen::trans randomization field");
			trn.print("Stimulus");
			mbox.put(trn);
			#5;
		end
		-> completed;
    endtask 

endclass //Sequencer






//////////////////////////////////////////////////////////////
////////////////         Driver Class          ///////////////
//////////////////////////////////////////////////////////////
class driver;

//    Resposible for driving transactions to the DUT through the virtual interface

	// Events that stops the write and read operations 
	event write_ended;
	event read_ended;
	
	
	// Creating virtual interface handle 
	virtual memory_if mem_vif;
	
	
	// Creating Mailbox handle
	mailbox mbox;

	// Transcations Counter 
	int trans_count;
	
	// Constructor 
	function new(virtual memory_if mem_vif, mailbox mbox);

		// Geting the interface 
		this.mem_vif = mem_vif;
		
		// Getting the mailbox handle from  environment 
		this.mbox = mbox;

	endfunction //new()

	// Adding a reset task, which initializes the Interface signals to default values
	task reset();
	
		wait(!mem_vif.Rst_n);
		
		$display("Time = %0t --------- Drivier Reset Task Started --------- \n", $time);
		
		`DRIV_IF.Wr_En   <= 'b0;
		`DRIV_IF.Rd_En   <= 'b0;
		`DRIV_IF.Data_in <= 'b0;
		`DRIV_IF.Address <= 'b0;
		
		wait(mem_vif.Rst_n);
		$display("Time = %0t --------- Drivier Reset Task Ended   --------- \n", $time);
			
	endtask


	// Driving the transaction items to the memory interface 
	task drive();
		
		$display("T = %0t [Driver] Starting .... \n", $time);
		forever
		begin

			Transaction #(32,5)trans;
			
			`DRIV_IF.Wr_En <= 'b0;
			`DRIV_IF.Rd_En <= 'b0;
			
			mbox.get(trans);
			
			$display("\n --- [Driver-Transfer: %0d] --- ", trans_count);
		
			@(posedge mem_vif.DRIVER.CLK);
				`DRIV_IF.Address <= trans.Address;

			// Write Operation 
			if(trans.Wr_En)
			begin
			
				`DRIV_IF.Wr_En 	 <= trans.Wr_En;
				`DRIV_IF.Data_in <= trans.Data_in;
				
				$display("Time = %0t --------------- Write Operation --------------- ",$time);
				$display("Wr_En = %0d \t Address = %0d \t Data_in = %0h",trans.Wr_En, trans.Address, trans.Data_in);
				
				@(posedge mem_vif.DRIVER.CLK);
			end
		

			// Read Operation 
			if(trans.Rd_En)
			begin

				`DRIV_IF.Rd_En <= trans.Rd_En;
				
				@(posedge mem_vif.DRIVER.CLK);
				`DRIV_IF.Rd_En <= 'b0;
				
				@(posedge mem_vif.DRIVER.CLK);
				trans.Data_out  <= `DRIV_IF.Data_out;
				trans.Valid_out <= `DRIV_IF.Valid_out;
				
				$display("Time = %0t --------------- Read Operation --------------- ",$time);
				$display("Rd_En = %0d \t Address = %0d \t Data_out = %0h \t Valid_out = %d",trans.Rd_En, `DRIV_IF.Address, `DRIV_IF.Data_out, `DRIV_IF.Valid_out);

			end
			trans_count++;
		end


	endtask 

endclass //driver





//////////////////////////////////////////////////////////////
////////////////         Monitor Class         ///////////////
//////////////////////////////////////////////////////////////
class Monitor;

/*

	** Samples the interface signals and converts the signal level activity to the transaction level
	** Send the sampled transaction to Scoreboard via Mailbox

*/


	// Virtual Memory Interface handle
	virtual memory_if mem_vif;
	
	
	
	// Mailbox from monitor into the subscriber
	mailbox mon_to_scb;
	
	
	
	// Constructor
	function new(virtual memory_if mem_vif, mailbox mon_to_scb);
	
		// Getting the Memory Interface
		this.mem_vif = mem_vif;
		
		// Getting the mailbox handles from the Environment Class
		this.mon_to_scb = mon_to_scb;
		
	endfunction
	
	
	
	
	// Sampling logic and sending the sampled transaction to the scoreboard
	task mont_task;
	
		forever
		begin
		
			Transaction #(32,5)trans;
			trans = new();
			
			
			@(posedge mem_vif.MONITOR.CLK)
			wait(`MONT_IF.Rd_En || `MONT_IF.Wr_En);
				
				trans.Wr_En   <= `MONT_IF.Wr_En;
				trans.Data_in <= `MONT_IF.Data_in;
				trans.Address <= `MONT_IF.Address;
				
				if(`MONT_IF.Rd_En)
				begin
				
					trans.Rd_En <= `MONT_IF.Rd_En;
					@(posedge mem_vif.MONITOR.CLK);
					@(posedge mem_vif.MONITOR.CLK);
					trans.Data_out  <= `MONT_IF.Data_out;
					trans.Valid_out <= `MONT_IF.Valid_out;
				
				end
		
			mon_to_scb.put(trans);
		end
	
	endtask

endclass





//////////////////////////////////////////////////////////////
////////////////       Scoreboard Class        ///////////////
//////////////////////////////////////////////////////////////
class Scoreboard;

/*
	
	Scoreboard receives the sampled packet from monitor,

		- if the transaction type is “read”, compares the read data with the local memory data
		- if the transaction type is “write”, local memory will be written with the wdata

*/


	// Mailbox handle
	mailbox mon_to_scb;
	
	
	// An integer to count the number of transactions
	int trans_count;
	

	// Creating an array that will be used as a local memory
	bit [31:0]loc_mem[31:0];
	
	
	function new(mailbox mon_to_scb);
	
		// Getting the mailbox handles from environment class
		this.mon_to_scb = mon_to_scb;
		
	endfunction
	
	
	
	// Storing wdata and compare rdata with stored data
	task scb_task;
	
	
		// Creating an instance of the Transaction Class
		Transaction #(32,5)trans;	
				
		forever
		begin
		
			#50;
			
			mon_to_scb.get(trans);
	
			if(trans.Wr_En)
			begin
			
				loc_mem[trans.Address] = trans.Data_in;
			
			end
			else if(trans.Rd_En)
			begin
				
				if(loc_mem[trans.Address] != trans.Data_out)
				$error("T = %0t, Sucsriber Failed: \nAddr = %d \nData :: Expected = %h \t Actual = %h", $time, trans.Address, loc_mem[trans.Address], trans.Data_out);
				else
				$display("Sucsriber Successeded !\n Addr = %0d Data :: Expected = %0h \t Actual = %0h", trans.Address, loc_mem[trans.Address], trans.Data_out);
			
			end


			trans_count++;
		
		end
	
	endtask
	
endclass





//////////////////////////////////////////////////////////////
////////////////       Environment Class       ///////////////
//////////////////////////////////////////////////////////////
class environment;

/*
	It is a container class, contains Mailbox, Sequencer, and Driver calsses

*/


	// Sequencer, Driver, Monitor and Subscriber Instances 
	Sequencer  Seq ;
	driver 	   drv ;
	Monitor    mont;
	Scoreboard scb ;
	

	
	// Virtual interface 
	virtual memory_if mem_vif;
	
	// Mailbox handle
	mailbox mbox;
	mailbox mon_to_scb;
	
	
	// Synchronize between the Drvier and the Sequencer through an Event
	event sync;
	
	
	function new(virtual memory_if mem_vif );
	
		// Get the interface from the test
		this.mem_vif = mem_vif;
		
		// Creating a mailbox handle, it will be shared across the Sequencer and Driver
		mbox = new();
		mon_to_scb = new();
		
		
		// Creating the Sequencer, Driver, Monitor, and Scoreboard
		Seq  = new(mbox, sync);
		drv  = new(mem_vif, mbox);
		mont = new(mem_vif, mon_to_scb);
		scb  = new(mon_to_scb);
		
	endfunction

	/*
	
		For better accessibility: I will divide the test operation on 3 tasks
		
		1. pre-test  task --> Method to call the initialization reset task
		2. test      task --> Method to generate the stimulus and drive it to the memory interface 
		3. post-test task --> Method to wait for the compeletion of the Sequencer and Driver operations 
	
	*/
	
	task pre_test();
	
		drv.reset();
	
	endtask
		
	
	task test;
	
		fork
		
			Seq.stimulus();
			drv.drive();
			mont.mont_task();
			scb.scb_task();
		
		join_any
		
	endtask
	
	
	task post_test;
	
		wait(sync.triggered);
		wait(Seq.repeat_count == drv.trans_count);
		wait(Seq.repeat_count == scb.trans_count);
		
	endtask


	// Test Run Task 
	task run();
	
		pre_test();
		test();
		post_test();
		
		$finish;
	
	endtask
	
endclass




//////////////////////////////////////////////////////////////
////////////////         Test Program          ///////////////
//////////////////////////////////////////////////////////////

// 1. Random Test 

program test(memory_if intf);

	class my_trans extends Transaction;
    
		bit [1:0] count;
		
		function void pre_randomize();
		  Wr_En.rand_mode(0);
		  Rd_En.rand_mode(0);
		  Address.rand_mode(0);
				
		  if(cnt %2 == 0) begin
			Wr_En = 1;
			Rd_En = 0;
			Address  = count;      
		  end 
		  else begin
			Wr_En = 0;
			Rd_En = 1;
			Address  = count;
			count++;
		  end
		  cnt++;
		endfunction
    
    endclass
	
	// Environment Class instance 
	environment env;
	my_trans    tr;
	
	initial
	begin
	
		// Environment Class handle Creation
		env = new(intf);
	
		tr = new();
		
		// Setting number of needed packets
		env.Seq.repeat_count = 50;				// Generate 15 packets
	
		// Calling the run test task from the Environment Class
		env.run();
		
	end
	
	
	
endprogram


/*
// 2. Write Read Test

	// postrandomize function, displaying randomized values of items 
	function void post_randomize();
		$display("--------- [Trans] post_randomize ------");
		if(Wr_En) $display("\t Address  = %0d\t wr_en = %d\t Data_in = %d",Address,Wr_En,Data_in);
		if(Rd_En) $display("\t Address  = %0h\t Rd_En = %d",Address,Rd_En);
		$display("-----------------------------------------");
	endfunction 
	
program test(mem_intf intf);
  
  class my_trans extends Transaction;
    
    bit [1:0] count;
    
    function void pre_randomize();
      Wr_En.rand_mode(0);
      Rd_En.rand_mode(0);
      Address.rand_mode(0);
            
      if(cnt %2 == 0) begin
        Wr_En = 1;
        Rd_En = 0;
        Address  = count;      
      end 
      else begin
        Wr_En = 0;
        Rd_En = 1;
        Address  = count;
        count++;
      end
      cnt++;
    endfunction
    
  endclass
    
  //declaring environment instance
  environment env;
  my_trans my_tr;
  
  initial begin
    //creating environment
    env = new(intf);
    
    my_tr = new();
    
    //setting the repeat count of generator as 4, means to generate 4 packets
    env.drv.repeat_count = 10;
    
    env.drv.trans = my_tr;
    
    //calling run of env, it interns calls generator and driver main tasks.
    env.run();
  end
endprogram
*/
